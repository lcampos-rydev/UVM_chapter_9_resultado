package gpio_agent_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

 
  `include "gpio_seq_item.svh"
  `include "gpio_driver.svh"
  `include "gpio_monitor.svh"
  `include "gpio_agent.svh"
  

endpackage